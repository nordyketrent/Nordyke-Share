//==============================================================================================================================================================
// grey_code
// Convert binary code to grey code
//
//  binary     grey
//   0000      0000
//   0001      0001
//   0010      0011
//   0011      0010
//   0100      0110
//   0101      0111
//   0110      0101
//   0111      0100
//   1000      1000
//   1001      1001
//   1010      1011
//   1011      1010
//   1100      1110
//   1101      1111
//   1110      1101
//   1111      1100
// 
//==============================================================================================================================================================

module grey_code #( parameter SIZE = 3 )
(
 input  [SIZE-1:0] binary_in,
 output [SIZE-1:0] grey_out
);

assign grey_out[SIZE-1:0] = binary_in[SIZE-1:0] ^ {1'b0,binary_in[SIZE-1:1]};

endmodule





